package sound_pkg;

    localparam int SOUND_ADDR [0:24] = '{
        20'd40000, // 音效0地址
        20'd120000, // 音效1地址
        20'h00000,  // 音效2地址
        20'd160000,  // 音效3地址
        20'h00000,  // 音效4地址
        20'd80000,  // 音效5地址
        20'd0,  // 音效6地址
        20'h00000,  // 音效7地址
        20'd200000,  // 音效8地址
        20'h00000,  // 音效9地址
        20'h00000,  // 音效10地址
        20'h00000,  // 音效11地址
        20'h00000,  // 音效12地址
        20'h00000,  // 音效13地址
        20'h00000,  // 音效14地址
        20'h00000,  // 音效15地址
        20'h00000,  // 音效16地址
        20'h00000,  // 音效17地址
        20'h00000,  // 音效18地址
        20'h00000,  // 音效19地址
        20'h00000,  // 音效20地址
        20'h00000,  // 音效21地址
        20'h00000,  // 音效22地址
        20'h00000,  // 音效23地址
        20'h00000   // 音效24地址
    };

    localparam logic [19:0] SOUND_LENGTH [0:24] = '{
        20'd39000, // 音效0長度
        20'd39000,  // 音效1長度
        20'h00000, // 音效2長度
        20'd39000, // 音效3長度
        20'h00000, // 音效4長度
        20'd39000, // 音效5長度
        20'd39000, // 音效6長度
        20'h00000, // 音效7長度
        20'd38000, // 音效8長度
        20'h00000, // 音效9長度
        20'h00000, // 音效10長度
        20'h00000, // 音效11長度
        20'h00000, // 音效12長度
        20'h00000, // 音效13長度
        20'h00000, // 音效14長度
        20'h00000, // 音效15長度
        20'h00000, // 音效16長度
        20'h00000, // 音效17長度
        20'h00000, // 音效18長度
        20'h00000, // 音效19長度
        20'h00000, // 音效20長度
        20'h00000, // 音效21長度
        20'h00000, // 音效22長度
        20'h00000, // 音效23長度
        20'h00000  // 音效24長度
    };

endpackage


