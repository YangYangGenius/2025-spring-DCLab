moudule SineWave(
    input i_clk,
    input i_rst_n,
    output [15:0] sine_out
);

    

endmodule